package clk_pkg; //bottom -> up order
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "seq.sv"
`include "driver.sv"
`include "agent.sv"
`include "sequencer.sv"
`include "clk_env.sv"
`include "base_test.sv"
endpackage
